-- datapath_aubie.vhd

-- entity reg_file (lab 2)
use work.dlx_types.all;
use work.bv_arithmetic.all;

entity reg_file is
    generic(prop_delay : Time := 5 ns);
    port (
        data_in     :   in dlx_word;
        readnotwrite:   in bit;
        clock       :   in bit;
	data_out    :   out dlx_word;
        reg_number  :   in register_index
    );
end entity reg_file;

---------------------------------------------
-- BEGIN Defining ARCHITECTURE "reg_file"  --
---------------------------------------------
architecture behavior of reg_file is
		----------------------------------------------------------
		-- 	Type Define (Act as 'storage' for our process)  --
		-- reg_type: defines a data structure for		--
		--	         an array of 32-bit words 		--
		----------------------------------------------------------
		type reg_type is array (0 to 31) of dlx_word;
begin
	reg_file_process: process(readnotwrite, clock, reg_number, data_in) is
	----------------------------------------------------------------------
	-- NOTE: Process accepts only input signals from our defined entity --
	----------------------------------------------------------------------
		----------------------------------------------------------
		-- 	Variable (Act as 'storage' for our process)  	--
		-- registers: implements reg_type and initializes       --
		--	      registers we use for this process		--
		----------------------------------------------------------
		variable registers: reg_type;
	begin
		-- Start process
		if (clock = '1') then
			if (readnotwrite = '1') then
				---------------------------------------------------------------
				-- 	[Performing "READ" Operation (readnotwrite = '1')]   --
				-- Here, we simply ignore 'data_in' and copy value in 	     --
				-- registers at index --> reg_number to data_out port signal --
				---------------------------------------------------------------
				data_out <= registers(bv_to_integer(reg_number)) after prop_delay;
			else
				------------------------------------------------------
				-- 	[Performing "WRITE" Operation]		    --
				-- Value from 'data_in' is copied into registers at --
				-- register index --> 'reg_number'		    --
				------------------------------------------------------
				registers(bv_to_integer(reg_number)) := data_in;
				------------------------------------------------------
				-- NOTE: No prop_delay is applied because we don't  --
				--	want to delay variable assignments. 	    --
				------------------------------------------------------
			end if;
		end if;
	end process reg_file_process;
end architecture behavior;


-- entity alu (lab 3)
use work.dlx_types.all;
use work.bv_arithmetic.all;

entity alu is
    generic(prop_delay : Time := 5 ns);
    port(
        operand1  :   in dlx_word;
        operand2  :   in dlx_word;
        operation :   in alu_operation_code;
        result    :   out dlx_word;
        error     :   out error_code
    );
end entity alu;

-- alu_operation_code values
-- 0000 unsigned add
-- 0001 signed add
-- 0010 2's compl add
-- 0011 2's compl sub
-- 0100 2's compl mul
-- 0101 2's compl divide
-- 0110 logical and
-- 0111 bitwise and
-- 1000 logical or
-- 1001 bitwise or
-- 1010 logical not (op1)
-- 1011 bitwise not (op1)
-- 1101-1111 output all zeros

-- error code values
-- 0000 = no error
-- 0001 = overflow (too big positive)
-- 0010 = underflow (too small neagative)
-- 0011 = divide by zero

architecture behavior of ALU is
    -- Define any types here that will be used

begin
    alu_process: process(operand1, operand2, operation) is
          -- Declare any local variables here
          variable temp_result: dlx_word := x"00000000";
          variable logical_true: dlx_word := x"00000001";
          variable logical_false: dlx_word := x"00000000";
          variable overflow_flag_set: boolean;
          variable div_by_zero: boolean;
          variable op1_logical_status: bit; -- 0 means false; 1 means true
          variable op2_logical_status: bit; -- 0 means false; 1 means true

          begin
              error <= "0000"; -- Default value for port signal output error
              case(operation) is
                  when "0000" => -- UNSIGNED ADD
                      bv_addu(operand1, operand2, temp_result, overflow_flag_set);
                      if overflow_flag_set then
                          error <= "0001";
                      end if;
                      result <= temp_result;
                  when "0001" => -- UNSIGNED SUBTRACT
                      bv_subu(operand1, operand2, temp_result, overflow_flag_set);
                      if overflow_flag_set then
                          error <= "0010";
                          -- Unsigned subtract is only concerned with underflow
                      end if;
                      result <= temp_result;
                  when "0010" => -- TWO'S COMPLEMENT ADD
                      bv_add(operand1, operand2, temp_result, overflow_flag_set);
                      if overflow_flag_set then
                          -- IF (+A) + (+B) = -C
                          if (operand1(31) = '0') AND (operand2(31) = '0') then
                              if (temp_result(31) = '1') then
                                  error <= "0001"; -- overflow occurred
                              end if;
                          -- (-A) + (-B) = +C
                          elsif (operand1(31) = '1') AND (operand2(31) = '1') then
                              if (temp_result(31) = '0') then
                                  error <= "0010"; -- underflow occurred
                              end if;
                          end if;
                      end if;
                      result <= temp_result;
                  when "0011" => -- TWO'S COMPLEMENT SUBTRACT
                      bv_sub(operand1, operand2, temp_result, overflow_flag_set);
                      if overflow_flag_set then
                          -- IF (-A) - (+B) = +C
                          if (operand1(31) = '1') AND (operand2(31) = '0') then
                              if (temp_result(31) = '0') then
                                  error <= "0010"; -- underflow occurred
                              end if;
                          -- IF (+A) - (-B) = -C
                          elsif (operand1(31) = '0') AND (operand2(31) = '1') then
                              if (temp_result(31) = '1') then
                                  error <= "0001"; -- overflow occurred
                              end if;
                          end if;
                      end if;
                      result <= temp_result;
                  when "0100" => -- TWO'S COMPLEMENT MULTIPLY - (2 underflow Conditions + 2 overflow conditions)
                      bv_mult(operand1, operand2, temp_result, overflow_flag_set);
                      if overflow_flag_set then
                          if (operand1(31) = '1') AND (operand2(31) = '0') then -- (-A x +B) = +C
                              error <= "0010"; -- underflow
                          elsif (operand1(31) = '0') AND (operand2(31) = '1') then -- (+A x -B) = +C
                              error <= "0010"; -- underflow
                          else -- (+A x +B) = -C OR (-A x -B) = -C
                              error <= "0001"; -- overflow
                          end if;
                      end if;
                      result <= temp_result;
                  when "0101" => -- TWO'S COMPLEMENT DIVIDE
                  ----------------------------------------------------------------------------------------
                  -- The only way a two's complement divide can underflow is if you divide the most
                  -- negative value by -ve 1. Divide underflow occurs when the divisor is much smaller
                  -- than the dividend. The result is almost zero. Test with 80000000 / FFFFFFFF
                  -- (Quotient will be smaller than the dividend)
                  -- NOTE: For grading purposes, this condition will not be tested but must be implemented
                  -----------------------------------------------------------------------------------------
                      bv_div(operand1, operand2, temp_result, div_by_zero, overflow_flag_set);
                      if div_by_zero then
                          error <= "0011"; --
                      elsif overflow_flag_set then
                          error <= "0010"; -- only an underflow can occur with divide (see note above)
                      end if;
                      result <= temp_result;
                  when "0110" => -- PERFORM LOGICAL AND
                  ------------------------------------------------------------------------
                  -- For logical operations, anything resulting in a non-zero value is 1,
                  -- for true. Anything resulting in all zeroes is assigned 0, false.
                  -- Logical operation always results in true (1) or false (0).
                  ------------------------------------------------------------------------
                      op1_logical_status := '0'; -- Default logical status for operand1
                      op2_logical_status := '0'; -- Default logical status for operand2
                      -- check if operand1 is a non-zero value --
                      for i in 31 downto 0 loop
                          -- If non-zero value, operand1 is logical true;
                          if (operand1(i) = '1') then
                              op1_logical_status := '1';
                              exit;
                          end if;
                      end loop;
                      -- check if operand2 is a non-zero value
                      for i in 31 downto 0 loop
                          -- If non-zero value, operand2 is logical true;
                          if (operand2(i) = '1') then
                              op2_logical_status := '1';
                              exit;
                          end if;
                      end loop;
                      -- IF operand statuses result in --> '1' && '1' = '1'
                      if ((op1_logical_status AND op2_logical_status) = '1') then
                          result <= logical_true; -- The result is logical true x"00000001"
                      else
                          result <= logical_false; -- Else result is logical false  x"00000000"
                      end if;
                  when "0111" => -- PERFORM BITWISE AND
                      for i in 31 downto 0 loop
                          temp_result(i) := operand1(i) AND operand2(i);
                      end loop;
                      result <= temp_result;
                  when "1000" => -- PERFORM LOGICAL OR
                  ------------------------------------------------------------------------
                  -- For logical operations, anything resulting in a non-zero value is 1,
                  -- for true. Anything resulting in a zero is assigned 0, false.
                  -- Logical operation always results in true (1) or false (0).
                  ------------------------------------------------------------------------
                      op1_logical_status := '0'; -- Default logical status for operand 1
                      op2_logical_status := '0'; -- Default logical status for operand 2
                      -- check if operand1 is a non-zero value --
                      for i in 31 downto 0 loop
                          -- If non-zero value, operand1 is logical true;
                          if (operand1(i) = '1') then
                              op1_logical_status := '1';
                              exit;
                          end if;
                      end loop;
                      -- check if operand2 is a non-zero value
                      for i in 31 downto 0 loop
                          -- If non-zero value, operand2 is logical true;
                          if (operand2(i) = '1') then
                              op2_logical_status := '1';
                              exit;
                          end if;
                      end loop;
                      -- IF operand statuses result in --> ('1'||'1' OR '1'||'0' OR '0'||'1' ) = '1'
                      if ((op1_logical_status OR op2_logical_status) = '1') then
                          result <= logical_true; -- The result is logical true x"00000001"
                      else
                          result <= logical_false; -- Else result is logical false  x"00000000"
                      end if;
                  when "1001" => -- PERFORM BITWISE OR
                      for i in 31 downto 0 loop
                          temp_result(i) := operand1(i) OR operand2(i);
                      end loop;
                      result <= temp_result;
                  when "1010" => -- PERFORM LOGICAL NOT OF OPERAND1 (ignore operand2)
                      temp_result := logical_true; -- Initially assigned to true (i.e. 32'h00000001)
                      for i in 31 downto 0 loop
                          if (NOT operand1(i) = '0') then -- i.e. IF operand1 is non-zero
                              temp_result := logical_false; -- logical NOT resulted in false; Therefore, NOT(operand1) = false
                              exit;
                          end if;
                      end loop;
                      result <= temp_result;
                  when "1011" => -- PERFORM BITWISE NOT OF OPERAND1 (ignore operand2)
                      for i in 31 downto 0 loop
                          temp_result(i) := NOT operand1(i);
                      end loop;
                      result <= temp_result;
                  when "1100" => -- CHECK IF OPERAND1 is zero
                      temp_result := logical_false;
                      if (operand1 = x"00000000") then
                          temp_result := logical_true;
                      end if;
                      result <= temp_result;
                  when others => -- 1101 thru 1111 outputs all zeroes
                      result <= x"00000000";
              end case;
   end process alu_process;
end architecture behavior;

-- entity dlx_register (lab 3)
use work.dlx_types.all;

entity dlx_register is
    generic(prop_delay : Time := 5 ns);
    port(
        in_val  :   in dlx_word;
        clock   :   in bit;
        out_val :   out dlx_word
    );
end entity dlx_register;

---------------------------------------------
-- BEGIN Defining ARCHITECTURE "dlx_register"  --
---------------------------------------------
architecture behavior of dlx_register is

begin
	dlx_reg_process: process(in_val, clock) is
	----------------------------------------------------------------------
	-- NOTE: Process accepts only input signals from our defined entity --
	----------------------------------------------------------------------
	begin
		-- Start process
		if (clock = '1') then
			out_val <= in_val after prop_delay;
		end if;
	end process dlx_reg_process;
end architecture behavior;

-- entity pcplusone
use work.dlx_types.all;
use work.bv_arithmetic.all;

entity pcplusone is
	generic(prop_delay: Time := 5 ns);
	port (
        input : in dlx_word;
        clock : in bit;
        output: out dlx_word
    );
end entity pcplusone;

architecture behavior of pcplusone is
begin
    plusone: process(input, clock) is  -- add clock input to make it execute
        variable newpc: dlx_word;
        variable error: boolean;
    begin
        if clock'event and clock = '1' then
            bv_addu(input,"00000000000000000000000000000001",newpc,error);
            output <= newpc after prop_delay;
        end if;
    end process plusone;
end architecture behavior;


-- entity mux
use work.dlx_types.all;

entity mux is
     generic(prop_delay : Time := 5 ns);
     port (
            input_1 : in dlx_word;
            input_0 : in dlx_word;
            which   : in bit;
            output  : out dlx_word
     );
end entity mux;

architecture behavior of mux is
begin
   muxProcess : process(input_1, input_0, which) is
   begin
      if (which = '1') then
         output <= input_1 after prop_delay;
      else
         output <= input_0 after prop_delay;
      end if;
   end process muxProcess;
end architecture behavior;
-- end entity mux

-- entity threeway_mux
use work.dlx_types.all;

entity threeway_mux is
    generic(prop_delay : Time := 5 ns);
    port (
        input_2 : in dlx_word;
        input_1 : in dlx_word;
        input_0 : in dlx_word;
        which   : in threeway_muxcode;
        output  : out dlx_word
    );
end entity threeway_mux;

architecture behavior of threeway_mux is
begin
   muxProcess : process(input_1, input_0, which) is
   begin
      if (which = "10" or which = "11" ) then
         output <= input_2 after prop_delay;
      elsif (which = "01") then
         output <= input_1 after prop_delay;
      else
         output <= input_0 after prop_delay;
      end if;
   end process muxProcess;
end architecture behavior;
-- end entity mux


-- entity memory
use work.dlx_types.all;
use work.bv_arithmetic.all;

entity memory is
    port (
        address       :   in dlx_word;
        readnotwrite  :   in bit;
        data_out      :   out dlx_word;
        data_in       :   in dlx_word;
        clock         :   in bit
    );
end memory;

architecture behavior of memory is

begin  -- behavior

    mem_behav: process(address,clock) is
    -- note that there is storage only for the first 1k of the memory, to speed
    -- up the simulation
        type memtype is array (0 to 1024) of dlx_word;
        variable data_memory : memtype;
    begin
    -- fill this in by hand to put some values in there
    -- some instructions
        data_memory(0) :=  X"30200000"; --LD R4, 0x100 -- [0011 0000 == x"30"] [0010 0 = x"4"][000 0000 0000 0000 0000]
        data_memory(1) :=  X"00000100"; -- address 0x100 for previous instruction

        data_memory(2) :=  X"30080000"; -- LD R1, 0x101
        data_memory(3) :=  X"00000101"; -- address 0x101 for previous instruction

        
        data_memory(4) :=  X"30100000"; -- LD R2, 0x102
        data_memory(5) :=  X"00000102"; -- address 0x102 for previous instruction

        -- This was initally data_memory(2) but I changed it to mem-address 6 so we can load R1 and R2 first
        data_memory(6) :=  "00000000000110000100010000000000"; -- ADDU R3,R1,R2

        -- note that this code runs every time an input signal to memory changes,
        -- so for testing, write to some other locations besides these
        data_memory(256) := "01010101000000001111111100000000";
        data_memory(257) := "10101010000000001111111100000000";
        data_memory(258) := "00000000000000000000000000000001";

                -- data_memory(259) - data_memory(1024) --


        if clock = '1' then
          if readnotwrite = '1' then
            -- do a read
            data_out <= data_memory(bv_to_natural(address)) after 5 ns;
          else
            -- do a write
            data_memory(bv_to_natural(address)) := data_in;
          end if;
        end if;
  end process mem_behav;
end behavior;
-- end entity memory
